module mips_reg_holder(
    input logic[31:0] reg_val_d,
    output logic[31:0] reg_val_q
);

endmodule


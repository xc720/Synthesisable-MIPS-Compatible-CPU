module mips_memory_data_register (
    input logic[31:0] memory_in,
    output logic[31:0] memory_out
) ;

endmodule

module mips_reg_holder(
    input logic[31:0] reg_val_d,
    output logic[31:0] reg_val_q
);

endmodule


module pc(
    input logic[31:0] pc_in,
    input logic pc_write_cond,
    input logic pc_write,
    input logic alu_zero,
    output logic[31:0] pc_out
);
    
endmodule
module pc(
    input logic[31:0] pc_in,
    output logic[31:0] pc_out
);


    assign pc_out = pc_in ;
    
endmodule
module mips_alu(
    input logic[31:0] a,
    input logic[31:0] b,
    output logic zero,
    output logic[31:0] alu_result
);

endmodule
